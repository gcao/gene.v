module gene

pub fn parse() {

}
