module types

pub struct Gene {
}