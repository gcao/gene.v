module gene

pub struct Parser {
	input str
}

(p &Parser) fn parse() {

}
